/*====================================
File name: seqinterfaceuence.sv
Date created: 18 March 2025
Description: interface component
====================================*/

interface our_interface(input logic clk);

    logic [7:0] input_1;
    logic [7:0] input_2;

    logic [15:0] output_3;
endinterface