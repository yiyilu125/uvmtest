/*====================================
File name: seqinterfaceuence.sv
Date created: 18 March 2025
Description: interface component
====================================*/

interface our_interface();

    //input_1
    //input_2
    
    //output_1
endinterface